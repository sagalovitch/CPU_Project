`timescale 1ns/10ps

module div32 (
    input wire [31:0] A,   // Dividend 
    input wire [31:0] M,   // Divisor 
    output reg [31:0] Q,   // Quotient 
    output reg [31:0] R    // Remainder 
);

    reg [63:0] temp;  
    integer i;  

    always @(*) begin
        Q = 0;
        temp = {32'b0, A};  

        if (M == 0) begin
            Q = 32'hFFFFFFFF;  
            R = 32'hFFFFFFFF;
        end else begin
            for (i = 0; i < 32; i = i + 1) begin
                temp = temp << 1;

                temp[63:32] = temp[63:32] - M;

                if (temp[63] == 1) begin

                    temp[63:32] = temp[63:32] + M;
                    Q = Q << 1;  
                end else begin
                    Q = (Q << 1) | 1; 
                end
            end
            R = temp[63:32];
        end
    end

endmodule
